../bios/bios.vh